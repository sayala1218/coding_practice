
module alwaysif2 (
    input      cpu_overheated,
    output reg shut_off_computer,
    input      arrived,
    input      gas_tank_empty,
    output reg keep_driving  ); //

    always_comb begin
        if (cpu_overheated)
           shut_off_computer = 1;
        else 
            shut_off_computer = 0;
    end

    always_comb begin
        if (~arrived)
           keep_driving = ~gas_tank_empty;
        else   
            keep_driving = ~arrived & ~gas_tank_empty;
    end

endmodule

// // synthesis verilog_input_version verilog_2001
// module alwyasif2 (
//     input      cpu_overheated,
//     output reg shut_off_computer,
//     input      arrived,
//     input      gas_tank_empty,
//     output reg keep_driving  ); //

//     always @(*) begin
//         if (cpu_overheated)
//            shut_off_computer = 1;
//         else 
//             shut_off_computer = 0;
//     end

//     always @(*) begin
//         if (~arrived)
//            keep_driving = ~gas_tank_empty;
//         else   
//             keep_driving = ~arrived & ~gas_tank_empty;
//     end

// endmodule